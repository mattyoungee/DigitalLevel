entity angleCalc is
port(

);

architecture logic of angleCalc is

end logic;