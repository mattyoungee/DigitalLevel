entity LEDcontrol is
port(

);

architecture logic of LEDcontrol is

end logic;